`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.07.2020 10:39:06
// Design Name: 
// Module Name: CLRX_wrapper
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CLRX_wrapper(

input        sys_clk,
input        RST_100_mb,
input        ap_rst_n,
input        rst,
input        rst_x,
input        rst_y,
input        rst_z,
input        clk_idelay_ref,
input        clk_x_p,
input        clk_y_p,
input        clk_z_p,
input        clk_x_n,
input        clk_y_n,
input        clk_z_n,
input [3:0]  serial_x_p, 
input [3:0]  serial_y_p, 
input [3:0]  serial_z_p, 
input [3:0]  serial_x_n, 
input [3:0]  serial_y_n, 
input [3:0]  serial_z_n,
input        LOCKED_x,
input        LOCKED_y,
input        LOCKED_z,
input        px_clk_x,
input        px_clk_y,
input        px_clk_z,
input        div2_clk_x,
input        div2_clk_y,
input        div2_clk_z,
input        div8_clk_x,
input        div8_clk_y,
input        div8_clk_z,
output       clk_x,
output       clk_y,
output       clk_z,
output       single_end_clk_x,
output       single_end_clk_y,
output       single_end_clk_z,
output [7:0] Ax,
output [7:0] Bx,
output [7:0] Cx,
output [7:0] Dy,
output [7:0] Ey,
output [7:0] Fy,
output [7:0] Gz,
output [7:0] Hz,
output [7:0] Iz,
output [3:0] LFDSx,
output [3:0] LFDSy,
output [3:0] LFDSz,
output       strb_ABC_val_x,
output       strb_DEF_val_y,
output       strb_GHI_val_z,
output       SOF_x,
output       SOF_dual_y,
output       EOL_x,
output       EOL_dual_y,
output [31:0] dna_high,
output [31:0] dna_low,
output        en_soc,
output [31:0] fifo_rst,
output [27:0] DATA_OUT0,
output [27:0] DATA_OUT1,
output [27:0] DATA_OUT2,
output        data_validx,
output        data_validy,
output  [15:0]   x_pcnt,   
output  [15:0]   x_lcnt,
output  [15:0]   y_pcnt,   
output  [15:0]   y_lcnt,

input  [8:0]  S_AXI_GPIO_araddr,
output        S_AXI_GPIO_arready,
input         S_AXI_GPIO_arvalid,
input  [8:0]  S_AXI_GPIO_awaddr,
output        S_AXI_GPIO_awready,
input         S_AXI_GPIO_awvalid,
input         S_AXI_GPIO_bready,
output [1:0]  S_AXI_GPIO_bresp,
output        S_AXI_GPIO_bvalid,
output [31:0] S_AXI_GPIO_rdata,
input         S_AXI_GPIO_rready,
output [1:0]  S_AXI_GPIO_rresp,
output        S_AXI_GPIO_rvalid,
input [31:0]  S_AXI_GPIO_wdata,
output        S_AXI_GPIO_wready,
input [3:0]   S_AXI_GPIO_wstrb,
input         S_AXI_GPIO_wvalid

    );
    
   
CLRX_wrapper_enc  CLRX_wrapper_enc (

.sys_clk(sys_clk),
.RST_100_mb(RST_100_mb),
.ap_rst_n(ap_rst_n),
.rst(rst),
.rst_x(rst_x),
.rst_y(rst_y),
.rst_z(rst_z),
.clk_idelay_ref(clk_idelay_ref),
.clk_x_p(clk_x_p),
.clk_y_p(clk_y_p),
.clk_z_p(clk_z_p),
.clk_x_n(clk_x_n),
.clk_y_n(clk_y_n),
.clk_z_n(clk_z_n),
.serial_x_p(serial_x_p),
.serial_y_p(serial_y_p),
.serial_z_p(serial_z_p),
.serial_x_n(serial_x_n),
.serial_y_n(serial_y_n),
.serial_z_n(serial_z_n),
.LOCKED_x(LOCKED_x),
.LOCKED_y(LOCKED_y),
.LOCKED_z(LOCKED_z),
.px_clk_x(px_clk_x),
.px_clk_y(px_clk_y),
.px_clk_z(px_clk_z),
.div2_clk_x(div2_clk_x),
.div2_clk_y(div2_clk_y),
.div2_clk_z(div2_clk_z),
.div8_clk_x(div8_clk_x),
.div8_clk_y(div8_clk_y),
.div8_clk_z(div8_clk_z),
.clk_x(clk_x),
.clk_y(clk_y),
.clk_z(clk_z),
.single_end_clk_x(single_end_clk_x),
.single_end_clk_y(single_end_clk_y),
.single_end_clk_z(single_end_clk_z),
.Ax(Ax),
.Bx(Bx),
.Cx(Cx),
.Dy(Dy),
.Ey(Ey),
.Fy(Fy),
.Gz(Gz),
.Hz(Hz),
.Iz(Iz),
.LFDSx(LFDSx),
.LFDSy(LFDSy),
.LFDSz(LFDSz),
.strb_ABC_val_x(strb_ABC_val_x),
.strb_DEF_val_y(strb_DEF_val_y),
.strb_GHI_val_z(strb_GHI_val_z),
.SOF_x(SOF_x),
.SOF_dual_y(SOF_dual_y),
.EOL_x(EOL_x),
.EOL_dual_y(EOL_dual_y),
.dna_high(dna_high),
.dna_low(dna_low),
.en_soc(en_soc),
.fifo_rst(fifo_rst),
.DATA_OUT0(DATA_OUT0),
.DATA_OUT1(DATA_OUT1),
.DATA_OUT2(DATA_OUT2),
.data_validx(data_validx),
.data_validy(data_validy),
.x_pcnt(x_pcnt),
.x_lcnt(x_lcnt),
.y_pcnt(y_pcnt),
.y_lcnt(y_lcnt),
.S_AXI_GPIO_araddr(S_AXI_GPIO_araddr),
.S_AXI_GPIO_arready(S_AXI_GPIO_arready),
.S_AXI_GPIO_arvalid(S_AXI_GPIO_arvalid),
.S_AXI_GPIO_awaddr(S_AXI_GPIO_awaddr),
.S_AXI_GPIO_awready(S_AXI_GPIO_awready),
.S_AXI_GPIO_awvalid(S_AXI_GPIO_awvalid),
.S_AXI_GPIO_bready(S_AXI_GPIO_bready),
.S_AXI_GPIO_bresp(S_AXI_GPIO_bresp),
.S_AXI_GPIO_bvalid(S_AXI_GPIO_bvalid),
.S_AXI_GPIO_rdata(S_AXI_GPIO_rdata),
.S_AXI_GPIO_rready(S_AXI_GPIO_rready),
.S_AXI_GPIO_rresp(S_AXI_GPIO_rresp),
.S_AXI_GPIO_rvalid(S_AXI_GPIO_rvalid),
.S_AXI_GPIO_wdata(S_AXI_GPIO_wdata),
.S_AXI_GPIO_wready(S_AXI_GPIO_wready),
.S_AXI_GPIO_wstrb(S_AXI_GPIO_wstrb),
.S_AXI_GPIO_wvalid(S_AXI_GPIO_wvalid)
);

endmodule
